--------------------------------------------------------------------------------
-- Title         : 8-Bit Full Adder
-- Project       : VHDL Synthesis Overview
-------------------------------------------------------------------------------
-- File          : eightBitAdder.vhd


