--------------------------------------------------------------------------------
-- Title         : 8-Bit Register
-- Project       : VHDL Synthesis Overview
-------------------------------------------------------------------------------
-- File          : eightBitRegister.vhd
