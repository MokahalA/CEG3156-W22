--------------------------------------------------------------------------------
-- Title         : Instruction Memory Block (ROM)
-- Project       : VHDL Synthesis Overview
-------------------------------------------------------------------------------
-- File          : instructionMemory.vhd

